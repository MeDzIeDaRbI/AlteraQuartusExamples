---------------------------------------------
-- PROJECT       : 7 Segments Display
-- ARBI MED ZIED : medzied.arbi@supcom.tn
-- WIEM HEDHILI  : wiem.hedhili@supcom.tn
-- SYSTEL B      : 08/02/2016
-- SUPCOM
---------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
---------------------------------------------
entity test is
	port (
				clk : in std_logic;
				bcd : in std_logic_vector(3 downto 0); --BCD input
				segment7 : out std_logic_vector(6 downto 0) -- 7 bit decoded output.
			);
end test;
---------------------------------------------
architecture Behavioral of test is
	component addN is
		generic(N: INTEGER:=4);
			port( A, B : in STD_LOGIC_VECTOR(N-1 downto 0);
					S : out STD_LOGIC_VECTOR(N downto 0));
		end component;
	
	begin
		G1: adder1 PORT MAP (A,B,S);
		process (clk,bcd)
			BEGIN
				if (clk'event and clk='1') then
					case bcd is
						when A<=(0) and B<=(0)=> segment7 <="0000001"; -- '0'
						when "0001"=> segment7 <="1001111"; -- '1'
						when "0010"=> segment7 <="0010010"; -- '2'
						when "0011"=> segment7 <="0000110"; -- '3'
						when "0100"=> segment7 <="1001100"; -- '4'
						when "0101"=> segment7 <="0100100"; -- '5'
						when "0110"=> segment7 <="0100000"; -- '6'
						when "0111"=> segment7 <="0001111"; -- '7'
						when "1000"=> segment7 <="0000000"; -- '8'
						when "1001"=> segment7 <="0000100"; -- '9'
						--nothing is displayed when a number more than 9 is given as input.
						when others=> segment7 <="1111111";
					end case;
				end if;
		end process;
		
end Behavioral;
